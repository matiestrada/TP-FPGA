library verilog;
use verilog.vl_types.all;
entity prueba_posicionamiento_vlg_vec_tst is
end prueba_posicionamiento_vlg_vec_tst;
