-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Wed Nov 27 18:34:51 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY giro_final IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        orientacion : IN STD_LOGIC_VECTOR(0 TO 1) := "00";
        dir_min : IN STD_LOGIC_VECTOR(0 TO 1) := "00";
        c_casilla : IN STD_LOGIC := '0';
        fin_giro : IN STD_LOGIC := '0';
        FW : OUT STD_LOGIC;
        girar : OUT STD_LOGIC;
        izq_der : OUT STD_LOGIC
    );
END giro_final;

ARCHITECTURE BEHAVIOR OF giro_final IS
    TYPE type_fstate IS (Check,giro_i,giro_d,avanzo);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,orientacion,dir_min,c_casilla,fin_giro)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Check;
            FW <= '0';
            girar <= '0';
            izq_der <= '0';
        ELSE
            FW <= '0';
            girar <= '0';
            izq_der <= '0';
            CASE fstate IS
                WHEN Check =>
                    IF ((((((((((orientacion(0 TO 1) = "00") AND (dir_min(0 TO 1) = "11")) OR ((orientacion(0 TO 1) = "01") AND (dir_min(0 TO 1) = "00"))) OR ((orientacion(0 TO 1) = "10") AND (dir_min(0 TO 1) = "01"))) OR ((orientacion(0 TO 1) = "11") AND (dir_min(0 TO 1) = "10"))) OR ((orientacion(0 TO 1) = "00") AND (dir_min(0 TO 1) = "10"))) OR ((orientacion(0 TO 1) = "01") AND (dir_min(0 TO 1) = "11"))) OR ((orientacion(0 TO 1) = "10") AND (dir_min(0 TO 1) = "00"))) OR ((orientacion(0 TO 1) = "11") AND (dir_min(0 TO 1) = "01")))) THEN
                        reg_fstate <= giro_i;
                    ELSIF ((((((orientacion(0 TO 1) = "00") AND (dir_min(0 TO 1) = "01")) OR ((orientacion(0 TO 1) = "01") AND (dir_min(0 TO 1) = "10"))) OR ((orientacion(0 TO 1) = "10") AND (dir_min(0 TO 1) = "11"))) OR ((orientacion(0 TO 1) = "11") AND (dir_min(0 TO 1) = "00")))) THEN
                        reg_fstate <= giro_d;
                    ELSIF ((orientacion(0 TO 1) = dir_min(0 TO 1))) THEN
                        reg_fstate <= avanzo;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Check;
                    END IF;

                    izq_der <= '0';

                    FW <= '0';

                    girar <= '0';
                WHEN giro_i =>
                    IF ((fin_giro = '1')) THEN
                        reg_fstate <= Check;
                    ELSIF ((fin_giro = '0')) THEN
                        reg_fstate <= giro_i;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= giro_i;
                    END IF;

                    izq_der <= '1';

                    FW <= '0';

                    girar <= '1';
                WHEN giro_d =>
                    IF ((fin_giro = '1')) THEN
                        reg_fstate <= Check;
                    ELSIF ((fin_giro = '0')) THEN
                        reg_fstate <= giro_d;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= giro_d;
                    END IF;

                    izq_der <= '0';

                    FW <= '0';

                    girar <= '1';
                WHEN avanzo =>
                    IF ((c_casilla = '1')) THEN
                        reg_fstate <= Check;
                    ELSIF ((c_casilla = '0')) THEN
                        reg_fstate <= avanzo;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= avanzo;
                    END IF;

                    izq_der <= '0';

                    FW <= '1';

                    girar <= '0';
                WHEN OTHERS => 
                    FW <= 'X';
                    girar <= 'X';
                    izq_der <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
