library verilog;
use verilog.vl_types.all;
entity pruebaparedes_vlg_vec_tst is
end pruebaparedes_vlg_vec_tst;
