library verilog;
use verilog.vl_types.all;
entity main is
    port(
        ADC_DIN         : out    vl_logic;
        clk0            : in     vl_logic;
        areset          : in     vl_logic;
        ADC_DOUT        : in     vl_logic;
        ADC_SCLK        : out    vl_logic;
        ADC_CS_N        : out    vl_logic;
        M1I             : out    vl_logic;
        clockcito       : in     vl_logic;
        RESET_GRAL      : in     vl_logic;
        orientacion     : out    vl_logic_vector(1 downto 0);
        Sensor_Frente   : in     vl_logic;
        pos             : out    vl_logic_vector(0 to 3);
        c_casilla       : out    vl_logic;
        Sensor_Linea    : in     vl_logic;
        M0I             : out    vl_logic;
        M1D             : out    vl_logic;
        M0D             : out    vl_logic;
        veld            : out    vl_logic;
        veli            : out    vl_logic;
        CONTADORRR      : out    vl_logic;
        dir_min         : out    vl_logic_vector(1 downto 0);
        Dir_Min12       : out    vl_logic_vector(1 downto 0);
        Dir_Min13       : out    vl_logic_vector(1 downto 0);
        Dir_Min14       : out    vl_logic_vector(1 downto 0);
        Dir_Min15       : out    vl_logic_vector(1 downto 0);
        Dir_Min2        : out    vl_logic_vector(1 downto 0);
        Dir_Min3        : out    vl_logic_vector(1 downto 0);
        Dir_Min4        : out    vl_logic_vector(1 downto 0);
        Dir_Min5        : out    vl_logic_vector(1 downto 0);
        Dir_Min6        : out    vl_logic_vector(1 downto 0);
        Dir_Min7        : out    vl_logic_vector(1 downto 0);
        Dir_Min8        : out    vl_logic_vector(1 downto 0);
        Dir_Min9        : out    vl_logic_vector(1 downto 0);
        \Dir_Min_10_\   : out    vl_logic_vector(1 downto 0);
        \Dir_Min_11_\   : out    vl_logic_vector(1 downto 0);
        \Dir_Min_1_\    : out    vl_logic_vector(1 downto 0);
        LEDS            : out    vl_logic_vector(7 downto 0);
        Mi_Peso12       : out    vl_logic_vector(3 downto 0);
        Mi_Peso13       : out    vl_logic_vector(3 downto 0);
        Mi_Peso14       : out    vl_logic_vector(3 downto 0);
        Mi_Peso15       : out    vl_logic_vector(3 downto 0);
        Mi_Peso2        : out    vl_logic_vector(3 downto 0);
        Mi_Peso3        : out    vl_logic_vector(3 downto 0);
        Mi_Peso4        : out    vl_logic_vector(3 downto 0);
        Mi_Peso5        : out    vl_logic_vector(3 downto 0);
        Mi_Peso6        : out    vl_logic_vector(3 downto 0);
        Mi_Peso7        : out    vl_logic_vector(3 downto 0);
        Mi_Peso8        : out    vl_logic_vector(3 downto 0);
        Mi_Peso9        : out    vl_logic_vector(3 downto 0);
        \Mi_Peso_0_\    : out    vl_logic_vector(3 downto 0);
        \Mi_Peso_10_\   : out    vl_logic_vector(3 downto 0);
        \Mi_Peso_11_\   : out    vl_logic_vector(3 downto 0);
        \Mi_Peso_1_\    : out    vl_logic_vector(3 downto 0)
    );
end main;
