library verilog;
use verilog.vl_types.all;
entity comp_prueba_vlg_vec_tst is
end comp_prueba_vlg_vec_tst;
