-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Tue Nov 26 12:47:37 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY control_prueba IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        I : IN STD_LOGIC := '0';
        D : IN STD_LOGIC := '0';
        F : IN STD_LOGIC := '0';
        estoy_fw : IN STD_LOGIC := '0';
        giro : OUT STD_LOGIC;
        IZQ_DER : OUT STD_LOGIC;
        FORWARD : OUT STD_LOGIC
    );
END control_prueba;

ARCHITECTURE BEHAVIOR OF control_prueba IS
    TYPE type_fstate IS (FW,GIRO_IZQ,GIRO_DER);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,I,D,F,estoy_fw)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= FW;
            giro <= '0';
            IZQ_DER <= '0';
            FORWARD <= '0';
        ELSE
            giro <= '0';
            IZQ_DER <= '0';
            FORWARD <= '0';
            CASE fstate IS
                WHEN FW =>
                    IF ((F = '0')) THEN
                        reg_fstate <= FW;
                    ELSIF (((((F = '1') AND (D = '1')) AND (I = '0')) OR (((F = '1') AND (D = '1')) AND (I = '1')))) THEN
                        reg_fstate <= GIRO_IZQ;
                    ELSIF (((((F = '1') AND (I = '1')) AND (D = '0')) OR (((F = '1') AND (I = '0')) AND (D = '0')))) THEN
                        reg_fstate <= GIRO_DER;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= FW;
                    END IF;

                    FORWARD <= '1';

                    IZQ_DER <= '0';

                    giro <= '0';
                WHEN GIRO_IZQ =>
                    IF ((estoy_fw = '0')) THEN
                        reg_fstate <= GIRO_IZQ;
                    ELSIF ((estoy_fw = '1')) THEN
                        reg_fstate <= FW;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= GIRO_IZQ;
                    END IF;

                    FORWARD <= '0';

                    IZQ_DER <= '1';

                    giro <= '1';
                WHEN GIRO_DER =>
                    IF ((estoy_fw = '0')) THEN
                        reg_fstate <= GIRO_DER;
                    ELSIF ((estoy_fw = '1')) THEN
                        reg_fstate <= FW;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= GIRO_DER;
                    END IF;

                    FORWARD <= '0';

                    IZQ_DER <= '0';

                    giro <= '1';
                WHEN OTHERS => 
                    giro <= 'X';
                    IZQ_DER <= 'X';
                    FORWARD <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
