-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Wed Nov 13 21:03:21 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY subsistema_3 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        y : IN STD_LOGIC := '0';
        cambio : IN STD_LOGIC := '0';
        pos : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END subsistema_3;

ARCHITECTURE BEHAVIOR OF subsistema_3 IS
    TYPE type_fstate IS (S00,S01,S02,S03,S10,S11,S12,S13,S20,S21,S22,S23,S30,S31,S32,S33);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x,y,cambio)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= S33;
            pos <= "0000";
        ELSE
            pos <= "0000";
            CASE fstate IS
                WHEN S00 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S01;
                    ELSIF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S00;
                    END IF;

                    pos <= "0000";
                WHEN S01 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S02;
                    ELSIF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S11;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S00;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S01;
                    END IF;

                    pos <= "0001";
                WHEN S02 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S03;
                    ELSIF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S12;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S01;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S02;
                    END IF;

                    pos <= "0010";
                WHEN S03 =>
                    IF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S13;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S02;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S03;
                    END IF;

                    pos <= "0011";
                WHEN S10 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S11;
                    ELSIF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S20;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S00;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S10;
                    END IF;

                    pos <= "0100";
                WHEN S11 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S12;
                    ELSIF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S21;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S01;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S11;
                    END IF;

                    pos <= "0101";
                WHEN S12 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S13;
                    ELSIF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S22;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S02;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S11;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S12;
                    END IF;

                    pos <= "0110";
                WHEN S13 =>
                    IF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S23;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S03;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S12;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S13;
                    END IF;

                    pos <= "0111";
                WHEN S20 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S21;
                    ELSIF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S30;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S20;
                    END IF;

                    pos <= "1000";
                WHEN S21 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S22;
                    ELSIF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S31;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S11;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S20;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S21;
                    END IF;

                    pos <= "1001";
                WHEN S22 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S23;
                    ELSIF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S32;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S12;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S21;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S22;
                    END IF;

                    pos <= "1010";
                WHEN S23 =>
                    IF ((((x = '1') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S33;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S13;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S22;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S23;
                    END IF;

                    pos <= "1011";
                WHEN S30 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S31;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S20;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S30;
                    END IF;

                    pos <= "1100";
                WHEN S31 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S32;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S21;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S30;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S31;
                    END IF;

                    pos <= "1101";
                WHEN S32 =>
                    IF ((((x = '0') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S33;
                    ELSIF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S22;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S31;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S32;
                    END IF;

                    pos <= "1110";
                WHEN S33 =>
                    IF ((((x = '0') AND (y = '0')) AND (cambio = '1'))) THEN
                        reg_fstate <= S23;
                    ELSIF ((((x = '1') AND (y = '1')) AND (cambio = '1'))) THEN
                        reg_fstate <= S32;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S33;
                    END IF;

                    pos <= "1111";
                WHEN OTHERS => 
                    pos <= "XXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
