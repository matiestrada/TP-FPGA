library verilog;
use verilog.vl_types.all;
entity prueba_control_vlg_vec_tst is
end prueba_control_vlg_vec_tst;
