library verilog;
use verilog.vl_types.all;
entity pared_vlg_vec_tst is
end pared_vlg_vec_tst;
