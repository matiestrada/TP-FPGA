library verilog;
use verilog.vl_types.all;
entity prueba_floodfill_vlg_vec_tst is
end prueba_floodfill_vlg_vec_tst;
