-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Mon Nov 11 16:53:37 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY subsistema_1 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        FW : IN STD_LOGIC := '0';
        I : IN STD_LOGIC := '0';
        D : IN STD_LOGIC := '0';
        M1I : OUT STD_LOGIC;
        M0I : OUT STD_LOGIC;
        M1D : OUT STD_LOGIC;
        M0D : OUT STD_LOGIC
    );
END subsistema_1;

ARCHITECTURE BEHAVIOR OF subsistema_1 IS
    TYPE type_fstate IS (Idle,Centrado,Pared_Izq,Pared_der);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,FW,I,D)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Idle;
            M1I <= '0';
            M0I <= '0';
            M1D <= '0';
            M0D <= '0';
        ELSE
            M1I <= '0';
            M0I <= '0';
            M1D <= '0';
            M0D <= '0';
            CASE fstate IS
                WHEN Idle =>
                    IF ((FW = '0')) THEN
                        reg_fstate <= Idle;
                    ELSIF ((((FW = '1') AND (I = '0')) AND (D = '0'))) THEN
                        reg_fstate <= Centrado;
                    ELSIF ((((FW = '1') AND (I = '1')) AND (D = '0'))) THEN
                        reg_fstate <= Pared_Izq;
                    ELSIF ((((FW = '1') AND (I = '0')) AND (D = '1'))) THEN
                        reg_fstate <= Pared_der;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Idle;
                    END IF;

                    M1D <= '0';

                    M1I <= '0';

                    M0D <= '0';

                    M0I <= '0';
                WHEN Centrado =>
                    IF ((FW = '0')) THEN
                        reg_fstate <= Idle;
                    ELSIF ((((FW = '1') AND (I = '1')) AND (D = '1'))) THEN
                        reg_fstate <= Centrado;
                    ELSIF ((((FW = '1') AND (I = '1')) AND (D = '0'))) THEN
                        reg_fstate <= Pared_Izq;
                    ELSIF ((((FW = '1') AND (I = '0')) AND (D = '1'))) THEN
                        reg_fstate <= Pared_der;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Centrado;
                    END IF;

                    M1D <= '0';

                    M1I <= '0';

                    M0D <= '1';

                    M0I <= '1';
                WHEN Pared_Izq =>
                    IF ((FW = '0')) THEN
                        reg_fstate <= Idle;
                    ELSIF ((((FW = '1') AND (I = '0')) AND (D = '0'))) THEN
                        reg_fstate <= Centrado;
                    ELSIF (((FW = '1') AND (I = '1'))) THEN
                        reg_fstate <= Pared_Izq;
                    ELSIF ((((FW = '1') AND (I = '0')) AND (D = '1'))) THEN
                        reg_fstate <= Pared_der;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Pared_Izq;
                    END IF;

                    M1D <= '0';

                    M1I <= '0';

                    M0D <= '0';

                    M0I <= '1';
                WHEN Pared_der =>
                    IF ((FW = '0')) THEN
                        reg_fstate <= Idle;
                    ELSIF ((((FW = '1') AND (I = '0')) AND (D = '0'))) THEN
                        reg_fstate <= Centrado;
                    ELSIF ((((FW = '1') AND (I = '1')) AND (D = '0'))) THEN
                        reg_fstate <= Pared_Izq;
                    ELSIF (((FW = '1') AND (D = '1'))) THEN
                        reg_fstate <= Pared_der;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Pared_der;
                    END IF;

                    M1D <= '0';

                    M1I <= '0';

                    M0D <= '1';

                    M0I <= '0';
                WHEN OTHERS => 
                    M1I <= 'X';
                    M0I <= 'X';
                    M1D <= 'X';
                    M0D <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
