library verilog;
use verilog.vl_types.all;
entity delay_5000_vlg_check_tst is
    port(
        fin_contador    : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end delay_5000_vlg_check_tst;
