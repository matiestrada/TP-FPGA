-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Nov 29 19:57:51 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY subsistema_3 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        ori : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        pos : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END subsistema_3;

ARCHITECTURE BEHAVIOR OF subsistema_3 IS
    TYPE type_fstate IS (S0,S1,S2,S3,S4,S5,S6,S7,S8,S9,S10,S11,S12,S13,S14,S15);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= S15;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,ori)
    BEGIN
        pos <= "0000";
        CASE fstate IS
            WHEN S0 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S1;
                ELSIF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S4;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S0;
                END IF;

                pos <= "0000";
            WHEN S1 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S2;
                ELSIF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S5;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S0;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S1;
                END IF;

                pos <= "0001";
            WHEN S2 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S3;
                ELSIF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S6;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S2;
                END IF;

                pos <= "0010";
            WHEN S3 =>
                IF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S7;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S2;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S3;
                END IF;

                pos <= "0011";
            WHEN S4 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S5;
                ELSIF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S8;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S0;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S4;
                END IF;

                pos <= "0100";
            WHEN S5 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S6;
                ELSIF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S9;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S1;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S4;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S5;
                END IF;

                pos <= "0101";
            WHEN S6 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S7;
                ELSIF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S10;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S2;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S5;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S6;
                END IF;

                pos <= "0110";
            WHEN S7 =>
                IF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S11;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S3;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S6;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S7;
                END IF;

                pos <= "0111";
            WHEN S8 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S9;
                ELSIF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S12;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S4;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S8;
                END IF;

                pos <= "1000";
            WHEN S9 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S10;
                ELSIF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S13;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S5;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S8;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S9;
                END IF;

                pos <= "1001";
            WHEN S10 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S11;
                ELSIF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S14;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S6;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S9;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S10;
                END IF;

                pos <= "1010";
            WHEN S11 =>
                IF ((ori(1 DOWNTO 0) = "10")) THEN
                    reg_fstate <= S15;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S7;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S10;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S11;
                END IF;

                pos <= "1011";
            WHEN S12 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S13;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S8;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S12;
                END IF;

                pos <= "1100";
            WHEN S13 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S14;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S9;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S12;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S13;
                END IF;

                pos <= "1101";
            WHEN S14 =>
                IF ((ori(1 DOWNTO 0) = "01")) THEN
                    reg_fstate <= S15;
                ELSIF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S10;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S13;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S14;
                END IF;

                pos <= "1110";
            WHEN S15 =>
                IF ((ori(1 DOWNTO 0) = "00")) THEN
                    reg_fstate <= S11;
                ELSIF ((ori(1 DOWNTO 0) = "11")) THEN
                    reg_fstate <= S14;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= S15;
                END IF;

                pos <= "1111";
            WHEN OTHERS => 
                pos <= "XXXX";
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
