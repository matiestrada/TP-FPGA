library verilog;
use verilog.vl_types.all;
entity Block5_vlg_vec_tst is
end Block5_vlg_vec_tst;
