library verilog;
use verilog.vl_types.all;
entity conexioooon_vlg_vec_tst is
end conexioooon_vlg_vec_tst;
