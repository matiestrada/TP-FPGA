library verilog;
use verilog.vl_types.all;
entity floodfill_para_simular_vlg_vec_tst is
end floodfill_para_simular_vlg_vec_tst;
