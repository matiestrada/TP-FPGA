library verilog;
use verilog.vl_types.all;
entity prueba_giro_vlg_vec_tst is
end prueba_giro_vlg_vec_tst;
