-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Nov 22 20:42:28 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Sistema_De_Orientacion IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        INFO_GIRO : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        orientacion : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
    );
END Sistema_De_Orientacion;

ARCHITECTURE BEHAVIOR OF Sistema_De_Orientacion IS
    TYPE type_fstate IS (NORTE,SUR,ESTE,OESTE,NORTE_IDLE,SUR_IDLE,ESTE_IDLE,OESTE_IDLE);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,INFO_GIRO)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= NORTE;
            orientacion <= "00";
        ELSE
            orientacion <= "00";
            CASE fstate IS
                WHEN NORTE =>
                    IF ((INFO_GIRO(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= NORTE_IDLE;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= NORTE;
                    END IF;
                WHEN SUR =>
                    IF ((INFO_GIRO(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= SUR_IDLE;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= SUR;
                    END IF;
                WHEN ESTE =>
                    IF ((INFO_GIRO(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= ESTE_IDLE;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ESTE;
                    END IF;
                WHEN OESTE =>
                    IF ((INFO_GIRO(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= OESTE_IDLE;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= OESTE;
                    END IF;
                WHEN NORTE_IDLE =>
                    IF ((INFO_GIRO(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= NORTE_IDLE;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "11")) THEN
                        reg_fstate <= SUR;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= OESTE;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= ESTE;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= NORTE_IDLE;
                    END IF;

                    orientacion <= "00";
                WHEN SUR_IDLE =>
                    IF ((INFO_GIRO(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= SUR_IDLE;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "11")) THEN
                        reg_fstate <= NORTE;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= ESTE;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= OESTE;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= SUR_IDLE;
                    END IF;

                    orientacion <= "10";
                WHEN ESTE_IDLE =>
                    IF ((INFO_GIRO(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= ESTE_IDLE;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "11")) THEN
                        reg_fstate <= OESTE;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= NORTE;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= SUR;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ESTE_IDLE;
                    END IF;

                    orientacion <= "01";
                WHEN OESTE_IDLE =>
                    IF ((INFO_GIRO(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= OESTE_IDLE;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "11")) THEN
                        reg_fstate <= ESTE;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= SUR;
                    ELSIF ((INFO_GIRO(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= NORTE;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= OESTE_IDLE;
                    END IF;

                    orientacion <= "11";
                WHEN OTHERS => 
                    orientacion <= "XX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
