library verilog;
use verilog.vl_types.all;
entity prueba_comparador_dir_vlg_check_tst is
    port(
        dir_correcta7   : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end prueba_comparador_dir_vlg_check_tst;
