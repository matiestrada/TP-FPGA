library verilog;
use verilog.vl_types.all;
entity prueba_comparador_dir_vlg_vec_tst is
end prueba_comparador_dir_vlg_vec_tst;
