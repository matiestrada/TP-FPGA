library verilog;
use verilog.vl_types.all;
entity delay_5000_vlg_vec_tst is
end delay_5000_vlg_vec_tst;
