-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Nov 28 17:31:51 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM3 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        c_casilla : IN STD_LOGIC := '0';
        forward : OUT STD_LOGIC;
        girar : OUT STD_LOGIC;
        izq_der : OUT STD_LOGIC
    );
END SM3;

ARCHITECTURE BEHAVIOR OF SM3 IS
    TYPE type_fstate IS (FW,check);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,c_casilla)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= FW;
            forward <= '0';
            girar <= '0';
            izq_der <= '0';
        ELSE
            forward <= '0';
            girar <= '0';
            izq_der <= '0';
            CASE fstate IS
                WHEN FW =>
                    IF ((c_casilla = '0')) THEN
                        reg_fstate <= FW;
                    ELSIF ((c_casilla = '1')) THEN
                        reg_fstate <= check;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= FW;
                    END IF;

                    forward <= '1';

                    izq_der <= '0';

                    girar <= '0';
                WHEN check =>
                    IF ((c_casilla = '0')) THEN
                        reg_fstate <= check;
                    ELSIF ((c_casilla = '1')) THEN
                        reg_fstate <= FW;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= check;
                    END IF;

                    forward <= '1';

                    izq_der <= '0';

                    girar <= '0';
                WHEN OTHERS => 
                    forward <= 'X';
                    girar <= 'X';
                    izq_der <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
