library verilog;
use verilog.vl_types.all;
entity prueba_orientacion_vlg_vec_tst is
end prueba_orientacion_vlg_vec_tst;
