-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Nov 21 16:49:50 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Sistema_De_Control_Prueba IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Pared_Delante : IN STD_LOGIC := '0';
        Fin_Giro : IN STD_LOGIC := '0';
        pared_der : IN STD_LOGIC := '0';
        pared_izq : IN STD_LOGIC := '0';
        FW : OUT STD_LOGIC;
        Girar : OUT STD_LOGIC;
        Izq_Der : OUT STD_LOGIC;
        giro180 : OUT STD_LOGIC
    );
END Sistema_De_Control_Prueba;

ARCHITECTURE BEHAVIOR OF Sistema_De_Control_Prueba IS
    TYPE type_fstate IS (Derecho,Giro_I,Giro_D,Giro_180);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Pared_Delante,Fin_Giro,pared_der,pared_izq)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Derecho;
            FW <= '0';
            Girar <= '0';
            Izq_Der <= '0';
            giro180 <= '0';
        ELSE
            FW <= '0';
            Girar <= '0';
            Izq_Der <= '0';
            giro180 <= '0';
            CASE fstate IS
                WHEN Derecho =>
                    IF ((Pared_Delante = '0')) THEN
                        reg_fstate <= Derecho;
                    ELSIF (((Pared_Delante = '1') AND (pared_izq = '0'))) THEN
                        reg_fstate <= Giro_I;
                    ELSIF ((((Pared_Delante = '1') AND (pared_der = '0')) AND (pared_izq = '1'))) THEN
                        reg_fstate <= Giro_D;
                    ELSIF ((((Pared_Delante = '1') AND (pared_der = '1')) AND (pared_izq = '1'))) THEN
                        reg_fstate <= Giro_180;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Derecho;
                    END IF;

                    giro180 <= '0';

                    Girar <= '0';

                    Izq_Der <= '1';

                    FW <= '1';
                WHEN Giro_I =>
                    IF ((Fin_Giro = '0')) THEN
                        reg_fstate <= Giro_I;
                    ELSIF ((Fin_Giro = '1')) THEN
                        reg_fstate <= Derecho;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Giro_I;
                    END IF;

                    giro180 <= '0';

                    Girar <= '1';

                    Izq_Der <= '1';

                    FW <= '0';
                WHEN Giro_D =>
                    IF ((Fin_Giro = '0')) THEN
                        reg_fstate <= Giro_D;
                    ELSIF ((Fin_Giro = '1')) THEN
                        reg_fstate <= Derecho;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Giro_D;
                    END IF;

                    giro180 <= '0';

                    Girar <= '1';

                    Izq_Der <= '0';

                    FW <= '0';
                WHEN Giro_180 =>
                    IF ((Fin_Giro = '0')) THEN
                        reg_fstate <= Giro_180;
                    ELSIF ((Fin_Giro = '1')) THEN
                        reg_fstate <= Derecho;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Giro_180;
                    END IF;

                    giro180 <= '1';

                    Girar <= '1';

                    Izq_Der <= '1';

                    FW <= '0';
                WHEN OTHERS => 
                    FW <= 'X';
                    Girar <= 'X';
                    Izq_Der <= 'X';
                    giro180 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
