library verilog;
use verilog.vl_types.all;
entity contador_7600_vlg_check_tst is
    port(
        fin_contador    : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end contador_7600_vlg_check_tst;
