library verilog;
use verilog.vl_types.all;
entity main_vlg_check_tst is
    port(
        ADC_CS_N        : in     vl_logic;
        ADC_DIN         : in     vl_logic;
        ADC_SCLK        : in     vl_logic;
        c_casilla       : in     vl_logic;
        CONTADORRR      : in     vl_logic;
        dir_min         : in     vl_logic_vector(1 downto 0);
        Dir_Min2        : in     vl_logic_vector(1 downto 0);
        Dir_Min3        : in     vl_logic_vector(1 downto 0);
        Dir_Min4        : in     vl_logic_vector(1 downto 0);
        Dir_Min5        : in     vl_logic_vector(1 downto 0);
        Dir_Min6        : in     vl_logic_vector(1 downto 0);
        Dir_Min7        : in     vl_logic_vector(1 downto 0);
        Dir_Min8        : in     vl_logic_vector(1 downto 0);
        Dir_Min9        : in     vl_logic_vector(1 downto 0);
        Dir_Min12       : in     vl_logic_vector(1 downto 0);
        Dir_Min13       : in     vl_logic_vector(1 downto 0);
        Dir_Min14       : in     vl_logic_vector(1 downto 0);
        Dir_Min15       : in     vl_logic_vector(1 downto 0);
        \Dir_Min_1_\    : in     vl_logic_vector(1 downto 0);
        \Dir_Min_10_\   : in     vl_logic_vector(1 downto 0);
        \Dir_Min_11_\   : in     vl_logic_vector(1 downto 0);
        LEDS            : in     vl_logic_vector(7 downto 0);
        M0D             : in     vl_logic;
        M0I             : in     vl_logic;
        M1D             : in     vl_logic;
        M1I             : in     vl_logic;
        Mi_Peso2        : in     vl_logic_vector(3 downto 0);
        Mi_Peso3        : in     vl_logic_vector(3 downto 0);
        Mi_Peso4        : in     vl_logic_vector(3 downto 0);
        Mi_Peso5        : in     vl_logic_vector(3 downto 0);
        Mi_Peso6        : in     vl_logic_vector(3 downto 0);
        Mi_Peso7        : in     vl_logic_vector(3 downto 0);
        Mi_Peso8        : in     vl_logic_vector(3 downto 0);
        Mi_Peso9        : in     vl_logic_vector(3 downto 0);
        Mi_Peso12       : in     vl_logic_vector(3 downto 0);
        Mi_Peso13       : in     vl_logic_vector(3 downto 0);
        Mi_Peso14       : in     vl_logic_vector(3 downto 0);
        Mi_Peso15       : in     vl_logic_vector(3 downto 0);
        \Mi_Peso_0_\    : in     vl_logic_vector(3 downto 0);
        \Mi_Peso_1_\    : in     vl_logic_vector(3 downto 0);
        \Mi_Peso_10_\   : in     vl_logic_vector(3 downto 0);
        \Mi_Peso_11_\   : in     vl_logic_vector(3 downto 0);
        orientacion     : in     vl_logic_vector(1 downto 0);
        pos             : in     vl_logic_vector(0 to 3);
        veld            : in     vl_logic;
        veli            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end main_vlg_check_tst;
