library verilog;
use verilog.vl_types.all;
entity cte1 is
    port(
        CONST_OUT       : out    vl_logic_vector(3 downto 0)
    );
end cte1;
