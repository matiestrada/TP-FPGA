-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Nov 21 14:44:05 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Detector_Cambio_Casilla IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Negro : IN STD_LOGIC := '0';
        Hab_Detector : IN STD_LOGIC := '0';
        Fin_Cont : IN STD_LOGIC := '0';
        Cambie_Casilla : OUT STD_LOGIC;
        Inicio_Cont : OUT STD_LOGIC
    );
END Detector_Cambio_Casilla;

ARCHITECTURE BEHAVIOR OF Detector_Cambio_Casilla IS
    TYPE type_fstate IS (Idle,Detecto_Blanco,Detecto_Negro,Confirmo_N,Casilla_Cambiada);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Negro,Hab_Detector,Fin_Cont)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Idle;
            Cambie_Casilla <= '0';
            Inicio_Cont <= '0';
        ELSE
            Cambie_Casilla <= '0';
            Inicio_Cont <= '0';
            CASE fstate IS
                WHEN Idle =>
                    IF ((Hab_Detector = '0')) THEN
                        reg_fstate <= Idle;
                    ELSIF (((Hab_Detector = '1') AND (Negro = '0'))) THEN
                        reg_fstate <= Detecto_Blanco;
                    ELSIF (((Hab_Detector = '1') AND (Negro = '1'))) THEN
                        reg_fstate <= Detecto_Negro;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Idle;
                    END IF;

                    Cambie_Casilla <= '0';

                    Inicio_Cont <= '0';
                WHEN Detecto_Blanco =>
                    IF ((Negro = '1')) THEN
                        reg_fstate <= Detecto_Negro;
                    ELSIF ((Negro = '0')) THEN
                        reg_fstate <= Detecto_Blanco;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Detecto_Blanco;
                    END IF;

                    Cambie_Casilla <= '0';

                    Inicio_Cont <= '0';
                WHEN Detecto_Negro =>
                    IF (((Negro = '1') AND (Fin_Cont = '1'))) THEN
                        reg_fstate <= Confirmo_N;
                    ELSIF ((Negro = '0')) THEN
                        reg_fstate <= Detecto_Blanco;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Detecto_Negro;
                    END IF;

                    Cambie_Casilla <= '0';

                    Inicio_Cont <= '1';
                WHEN Confirmo_N =>
                    IF ((Negro = '1')) THEN
                        reg_fstate <= Confirmo_N;
                    ELSIF ((Negro = '0')) THEN
                        reg_fstate <= Casilla_Cambiada;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Confirmo_N;
                    END IF;

                    Cambie_Casilla <= '0';

                    Inicio_Cont <= '0';
                WHEN Casilla_Cambiada =>
                    reg_fstate <= Idle;

                    Cambie_Casilla <= '1';

                    Inicio_Cont <= '0';
                WHEN OTHERS => 
                    Cambie_Casilla <= 'X';
                    Inicio_Cont <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
