library verilog;
use verilog.vl_types.all;
entity Block5_vlg_check_tst is
    port(
        dir_correcta    : in     vl_logic;
        FW              : in     vl_logic;
        giro            : in     vl_logic;
        izq_der         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Block5_vlg_check_tst;
