-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Nov 29 00:14:04 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY control IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        dir_correcta : IN STD_LOGIC := '0';
        prioridad_i_d : IN STD_LOGIC := '0';
        fin_giro : IN STD_LOGIC := '0';
        pared_delante : IN STD_LOGIC := '0';
        FW : OUT STD_LOGIC;
        giro : OUT STD_LOGIC;
        izq_der : OUT STD_LOGIC
    );
END control;

ARCHITECTURE BEHAVIOR OF control IS
    TYPE type_fstate IS (check,giro_izq,giro_der,forward);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,dir_correcta,prioridad_i_d,fin_giro,pared_delante)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= check;
            FW <= '0';
            giro <= '0';
            izq_der <= '0';
        ELSE
            FW <= '0';
            giro <= '0';
            izq_der <= '0';
            CASE fstate IS
                WHEN check =>
                    IF (((dir_correcta = '0') AND (prioridad_i_d = '0'))) THEN
                        reg_fstate <= giro_izq;
                    ELSIF (((dir_correcta = '0') AND (prioridad_i_d = '1'))) THEN
                        reg_fstate <= giro_der;
                    ELSIF ((dir_correcta = '1')) THEN
                        reg_fstate <= forward;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= check;
                    END IF;

                    giro <= '0';

                    FW <= '0';

                    izq_der <= '0';
                WHEN giro_izq =>
                    IF ((fin_giro = '0')) THEN
                        reg_fstate <= giro_izq;
                    ELSIF ((fin_giro = '1')) THEN
                        reg_fstate <= check;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= giro_izq;
                    END IF;

                    giro <= '1';

                    FW <= '0';

                    izq_der <= '1';
                WHEN giro_der =>
                    IF ((fin_giro = '0')) THEN
                        reg_fstate <= giro_der;
                    ELSIF ((fin_giro = '1')) THEN
                        reg_fstate <= check;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= giro_der;
                    END IF;

                    giro <= '1';

                    FW <= '0';

                    izq_der <= '0';
                WHEN forward =>
                    IF (((dir_correcta = '1') AND (pared_delante = '0'))) THEN
                        reg_fstate <= forward;
                    ELSIF (((dir_correcta = '0') OR (pared_delante = '1'))) THEN
                        reg_fstate <= check;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= forward;
                    END IF;

                    giro <= '0';

                    FW <= '1';

                    izq_der <= '0';
                WHEN OTHERS => 
                    FW <= 'X';
                    giro <= 'X';
                    izq_der <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
