library verilog;
use verilog.vl_types.all;
entity contador_7600_vlg_vec_tst is
end contador_7600_vlg_vec_tst;
