library verilog;
use verilog.vl_types.all;
entity cte1_vlg_vec_tst is
end cte1_vlg_vec_tst;
