library verilog;
use verilog.vl_types.all;
entity contador_10_vlg_vec_tst is
end contador_10_vlg_vec_tst;
