library verilog;
use verilog.vl_types.all;
entity pRUEBAFF_vlg_vec_tst is
end pRUEBAFF_vlg_vec_tst;
